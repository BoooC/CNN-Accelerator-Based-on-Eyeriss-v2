// ====================================================================================================== //
// This module is router cluster.
// router cluster module inregrates 9 iact routers, 3 weight routers, 3 psum routers.
// This module is one of the main part in this accelerator architecture.
// Its iact   routers are connected to all PEs 			  in PE cluster (one-to-one). 
// Its weight routers are connected to all rows of PEs 	  in PE cluster (one-to-row). 
// Its psum   routers are connected to all columns of PEs in PE cluster (one=to-column). 
//
// router cluster is the core of Hierarchical mesh-NoC, which can provide flexibility to the accelerator.
// This architecture can support all types of data flow topology wiht data_in_sel and data_out_sel control signals.
// ====================================================================================================== //

module Router_Cluster(
	// ----------- control ----------- //
	input  [1:0]  iact_0_data_in_sel,
	input  [1:0]  iact_0_data_out_sel,
	input  [1:0]  iact_1_data_in_sel,
	input  [1:0]  iact_1_data_out_sel,
	input  [1:0]  iact_2_data_in_sel,
	input  [1:0]  iact_2_data_out_sel,
	
	input         weight_0_data_in_sel,
	input         weight_0_data_out_sel,
	input         weight_1_data_in_sel,
	input         weight_1_data_out_sel,
	input         weight_2_data_in_sel,
	input         weight_2_data_out_sel,
	
	input  		  psum_0_data_in_sel,
	input  		  psum_0_data_out_sel,
	input  		  psum_1_data_in_sel,
	input  		  psum_1_data_out_sel,
	input  		  psum_2_data_in_sel,
	input  		  psum_2_data_out_sel,
	
	// ----------- iact router 0_0 ----------- //
	// src port
	output        iact_0_0_GLB_address_in_ready,
	input         iact_0_0_GLB_address_in_valid,
	input  [6:0]  iact_0_0_GLB_address_in_bits,
	output        iact_0_0_GLB_data_in_ready,
	input         iact_0_0_GLB_data_in_valid,
	input  [11:0] iact_0_0_GLB_data_in_bits,
				
	output        iact_0_0_north_address_in_ready,
	input         iact_0_0_north_address_in_valid,
	input  [6:0]  iact_0_0_north_address_in_bits,
	output        iact_0_0_north_data_in_ready,
	input         iact_0_0_north_data_in_valid,
	input  [11:0] iact_0_0_north_data_in_bits,
					
	output        iact_0_0_south_address_in_ready,
	input         iact_0_0_south_address_in_valid,
	input  [6:0]  iact_0_0_south_address_in_bits,
	output        iact_0_0_south_data_in_ready,
	input         iact_0_0_south_data_in_valid,
	input  [11:0] iact_0_0_south_data_in_bits,
					
	output        iact_0_0_horiz_address_in_ready,
	input         iact_0_0_horiz_address_in_valid,
	input  [6:0]  iact_0_0_horiz_address_in_bits,
	output        iact_0_0_horiz_data_in_ready,
	input         iact_0_0_horiz_data_in_valid,                        
	input  [11:0] iact_0_0_horiz_data_in_bits,                          
	// dst port                                                    
	input         iact_0_0_PE_address_out_ready,                        
	output [6:0]  iact_0_0_PE_address_out_bits,                         
	output        iact_0_0_PE_address_out_valid,                        
	input         iact_0_0_PE_data_out_ready,
	output        iact_0_0_PE_data_out_valid,
	output [11:0] iact_0_0_PE_data_out_bits,
					
	input		  iact_0_0_north_address_out_ready,
	output        iact_0_0_north_address_out_valid,
	output [6:0]  iact_0_0_north_address_out_bits,
	input		  iact_0_0_north_data_out_ready,
	output        iact_0_0_north_data_out_valid,
	output [11:0] iact_0_0_north_data_out_bits,
				
	input         iact_0_0_south_address_out_ready, 
	output        iact_0_0_south_address_out_valid,  
	output [6:0]  iact_0_0_south_address_out_bits, 
	input         iact_0_0_south_data_out_ready,
	output        iact_0_0_south_data_out_valid,
	output [11:0] iact_0_0_south_data_out_bits,
					
	input         iact_0_0_horiz_address_out_ready, 
	output        iact_0_0_horiz_address_out_valid,  
	output [6:0]  iact_0_0_horiz_address_out_bits, 
	input         iact_0_0_horiz_data_out_ready,
	output        iact_0_0_horiz_data_out_valid,
	output [11:0] iact_0_0_horiz_data_out_bits,
	
	
	// ----------- iact router 0_1 ----------- //
	// src port
	output        iact_0_1_GLB_address_in_ready,
	input         iact_0_1_GLB_address_in_valid,
	input  [6:0]  iact_0_1_GLB_address_in_bits,
	output        iact_0_1_GLB_data_in_ready,
	input         iact_0_1_GLB_data_in_valid,
	input  [11:0] iact_0_1_GLB_data_in_bits,
						 
	output        iact_0_1_north_address_in_ready,
	input         iact_0_1_north_address_in_valid,
	input  [6:0]  iact_0_1_north_address_in_bits,
	output        iact_0_1_north_data_in_ready,
	input         iact_0_1_north_data_in_valid,
	input  [11:0] iact_0_1_north_data_in_bits,
						 
	output        iact_0_1_south_address_in_ready,
	input         iact_0_1_south_address_in_valid,
	input  [6:0]  iact_0_1_south_address_in_bits,
	output        iact_0_1_south_data_in_ready,
	input         iact_0_1_south_data_in_valid,
	input  [11:0] iact_0_1_south_data_in_bits,
						 
	output        iact_0_1_horiz_address_in_ready,
	input         iact_0_1_horiz_address_in_valid,
	input  [6:0]  iact_0_1_horiz_address_in_bits,
	output        iact_0_1_horiz_data_in_ready,
	input         iact_0_1_horiz_data_in_valid,                        
	input  [11:0] iact_0_1_horiz_data_in_bits,                          
	// dst port                                                      
	input         iact_0_1_PE_address_out_ready,                        
	output [6:0]  iact_0_1_PE_address_out_bits,                         
	output        iact_0_1_PE_address_out_valid,                        
	input         iact_0_1_PE_data_out_ready,
	output        iact_0_1_PE_data_out_valid,
	output [11:0] iact_0_1_PE_data_out_bits,
						 
	input		  iact_0_1_north_address_out_ready,
	output        iact_0_1_north_address_out_valid,
	output [6:0]  iact_0_1_north_address_out_bits,
	input		  iact_0_1_north_data_out_ready,
	output        iact_0_1_north_data_out_valid,
	output [11:0] iact_0_1_north_data_out_bits,
						 
	input         iact_0_1_south_address_out_ready, 
	output        iact_0_1_south_address_out_valid,  
	output [6:0]  iact_0_1_south_address_out_bits, 
	input         iact_0_1_south_data_out_ready,
	output        iact_0_1_south_data_out_valid,
	output [11:0] iact_0_1_south_data_out_bits,
						 
	input         iact_0_1_horiz_address_out_ready, 
	output        iact_0_1_horiz_address_out_valid,  
	output [6:0]  iact_0_1_horiz_address_out_bits, 
	input         iact_0_1_horiz_data_out_ready,
	output        iact_0_1_horiz_data_out_valid,
	output [11:0] iact_0_1_horiz_data_out_bits,
	
	
	// ----------- iact router 0_2 ----------- //
	// src port
	output        iact_0_2_GLB_address_in_ready,
	input         iact_0_2_GLB_address_in_valid,
	input  [6:0]  iact_0_2_GLB_address_in_bits,
	output        iact_0_2_GLB_data_in_ready,
	input         iact_0_2_GLB_data_in_valid,
	input  [11:0] iact_0_2_GLB_data_in_bits,
						 
	output        iact_0_2_north_address_in_ready,
	input         iact_0_2_north_address_in_valid,
	input  [6:0]  iact_0_2_north_address_in_bits,
	output        iact_0_2_north_data_in_ready,
	input         iact_0_2_north_data_in_valid,
	input  [11:0] iact_0_2_north_data_in_bits,
						 
	output        iact_0_2_south_address_in_ready,
	input         iact_0_2_south_address_in_valid,
	input  [6:0]  iact_0_2_south_address_in_bits,
	output        iact_0_2_south_data_in_ready,
	input         iact_0_2_south_data_in_valid,
	input  [11:0] iact_0_2_south_data_in_bits,
						
	output        iact_0_2_horiz_address_in_ready,
	input         iact_0_2_horiz_address_in_valid,
	input  [6:0]  iact_0_2_horiz_address_in_bits,
	output        iact_0_2_horiz_data_in_ready,
	input         iact_0_2_horiz_data_in_valid,                        
	input  [11:0] iact_0_2_horiz_data_in_bits,                          
	// dst port                                                    
	input         iact_0_2_PE_address_out_ready,                        
	output [6:0]  iact_0_2_PE_address_out_bits,                         
	output        iact_0_2_PE_address_out_valid,                        
	input         iact_0_2_PE_data_out_ready,
	output        iact_0_2_PE_data_out_valid,
	output [11:0] iact_0_2_PE_data_out_bits,
						 
	input		  iact_0_2_north_address_out_ready,
	output        iact_0_2_north_address_out_valid,
	output [6:0]  iact_0_2_north_address_out_bits,
	input		  iact_0_2_north_data_out_ready,
	output        iact_0_2_north_data_out_valid,
	output [11:0] iact_0_2_north_data_out_bits,
						 
	input         iact_0_2_south_address_out_ready, 
	output        iact_0_2_south_address_out_valid,  
	output [6:0]  iact_0_2_south_address_out_bits, 
	input         iact_0_2_south_data_out_ready,
	output        iact_0_2_south_data_out_valid,
	output [11:0] iact_0_2_south_data_out_bits,
						 
	input         iact_0_2_horiz_address_out_ready, 
	output        iact_0_2_horiz_address_out_valid,  
	output [6:0]  iact_0_2_horiz_address_out_bits, 
	input         iact_0_2_horiz_data_out_ready,
	output        iact_0_2_horiz_data_out_valid,
	output [11:0] iact_0_2_horiz_data_out_bits,
	
	
	// ----------- iact router 1_0 ----------- //
	// src port
	output        iact_1_0_GLB_address_in_ready,
	input         iact_1_0_GLB_address_in_valid,
	input  [6:0]  iact_1_0_GLB_address_in_bits,
	output        iact_1_0_GLB_data_in_ready,
	input         iact_1_0_GLB_data_in_valid,
	input  [11:0] iact_1_0_GLB_data_in_bits,
				
	output        iact_1_0_north_address_in_ready,
	input         iact_1_0_north_address_in_valid,
	input  [6:0]  iact_1_0_north_address_in_bits,
	output        iact_1_0_north_data_in_ready,
	input         iact_1_0_north_data_in_valid,
	input  [11:0] iact_1_0_north_data_in_bits,
					
	output        iact_1_0_south_address_in_ready,
	input         iact_1_0_south_address_in_valid,
	input  [6:0]  iact_1_0_south_address_in_bits,
	output        iact_1_0_south_data_in_ready,
	input         iact_1_0_south_data_in_valid,
	input  [11:0] iact_1_0_south_data_in_bits,
					
	output        iact_1_0_horiz_address_in_ready,
	input         iact_1_0_horiz_address_in_valid,
	input  [6:0]  iact_1_0_horiz_address_in_bits,
	output        iact_1_0_horiz_data_in_ready,
	input         iact_1_0_horiz_data_in_valid,         
	input  [11:0] iact_1_0_horiz_data_in_bits,          
	// dst port          0_                                            
	input         iact_1_0_PE_address_out_ready,        
	output        iact_1_0_PE_address_out_valid,         
	output [6:0]  iact_1_0_PE_address_out_bits,        
	input         iact_1_0_PE_data_out_ready,
	output        iact_1_0_PE_data_out_valid,
	output [11:0] iact_1_0_PE_data_out_bits,
					
	input		  iact_1_0_north_address_out_ready,
	output        iact_1_0_north_address_out_valid,
	output [6:0]  iact_1_0_north_address_out_bits,
	input		  iact_1_0_north_data_out_ready,
	output        iact_1_0_north_data_out_valid,
	output [11:0] iact_1_0_north_data_out_bits,
						
	input         iact_1_0_south_address_out_ready, 
	output        iact_1_0_south_address_out_valid,  
	output [6:0]  iact_1_0_south_address_out_bits, 
	input         iact_1_0_south_data_out_ready,
	output        iact_1_0_south_data_out_valid,
	output [11:0] iact_1_0_south_data_out_bits,
					
	input         iact_1_0_horiz_address_out_ready, 
	output        iact_1_0_horiz_address_out_valid,  
	output [6:0]  iact_1_0_horiz_address_out_bits, 
	input         iact_1_0_horiz_data_out_ready,
	output        iact_1_0_horiz_data_out_valid,
	output [11:0] iact_1_0_horiz_data_out_bits,
	
	
	// ----------- iact router 1_1 ----------- //
	// src port
	output        iact_1_1_GLB_address_in_ready,
	input         iact_1_1_GLB_address_in_valid,
	input  [6:0]  iact_1_1_GLB_address_in_bits,
	output        iact_1_1_GLB_data_in_ready,
	input         iact_1_1_GLB_data_in_valid,
	input  [11:0] iact_1_1_GLB_data_in_bits,
						 
	output        iact_1_1_north_address_in_ready,
	input         iact_1_1_north_address_in_valid,
	input  [6:0]  iact_1_1_north_address_in_bits,
	output        iact_1_1_north_data_in_ready,
	input         iact_1_1_north_data_in_valid,
	input  [11:0] iact_1_1_north_data_in_bits,
						 
	output        iact_1_1_south_address_in_ready,
	input         iact_1_1_south_address_in_valid,
	input  [6:0]  iact_1_1_south_address_in_bits,
	output        iact_1_1_south_data_in_ready,
	input         iact_1_1_south_data_in_valid,
	input  [11:0] iact_1_1_south_data_in_bits,
						 
	output        iact_1_1_horiz_address_in_ready,
	input         iact_1_1_horiz_address_in_valid,
	input  [6:0]  iact_1_1_horiz_address_in_bits,
	output        iact_1_1_horiz_data_in_ready,
	input         iact_1_1_horiz_data_in_valid,         
	input  [11:0] iact_1_1_horiz_data_in_bits,          
	// dst port                                                     
	input         iact_1_1_PE_address_out_ready,        
	output        iact_1_1_PE_address_out_valid,         
	output [6:0]  iact_1_1_PE_address_out_bits,        
	input         iact_1_1_PE_data_out_ready,
	output        iact_1_1_PE_data_out_valid,
	output [11:0] iact_1_1_PE_data_out_bits,
						 
	input		  iact_1_1_north_address_out_ready,
	output        iact_1_1_north_address_out_valid,
	output [6:0]  iact_1_1_north_address_out_bits,
	input		  iact_1_1_north_data_out_ready,
	output        iact_1_1_north_data_out_valid,
	output [11:0] iact_1_1_north_data_out_bits,
						 
	input         iact_1_1_south_address_out_ready, 
	output        iact_1_1_south_address_out_valid,  
	output [6:0]  iact_1_1_south_address_out_bits, 
	input         iact_1_1_south_data_out_ready,
	output        iact_1_1_south_data_out_valid,
	output [11:0] iact_1_1_south_data_out_bits,
						 
	input         iact_1_1_horiz_address_out_ready, 
	output        iact_1_1_horiz_address_out_valid,  
	output [6:0]  iact_1_1_horiz_address_out_bits, 
	input         iact_1_1_horiz_data_out_ready,
	output        iact_1_1_horiz_data_out_valid,
	output [11:0] iact_1_1_horiz_data_out_bits,
	
	
	// ----------- iact router 1_2 ----------- //
	// src port
	output        iact_1_2_GLB_address_in_ready,
	input         iact_1_2_GLB_address_in_valid,
	input  [6:0]  iact_1_2_GLB_address_in_bits,
	output        iact_1_2_GLB_data_in_ready,
	input         iact_1_2_GLB_data_in_valid,
	input  [11:0] iact_1_2_GLB_data_in_bits,
						 
	output        iact_1_2_north_address_in_ready,
	input         iact_1_2_north_address_in_valid,
	input  [6:0]  iact_1_2_north_address_in_bits,
	output        iact_1_2_north_data_in_ready,
	input         iact_1_2_north_data_in_valid,
	input  [11:0] iact_1_2_north_data_in_bits,
						 
	output        iact_1_2_south_address_in_ready,
	input         iact_1_2_south_address_in_valid,
	input  [6:0]  iact_1_2_south_address_in_bits,
	output        iact_1_2_south_data_in_ready,
	input         iact_1_2_south_data_in_valid,
	input  [11:0] iact_1_2_south_data_in_bits,
						 
	output        iact_1_2_horiz_address_in_ready,
	input         iact_1_2_horiz_address_in_valid,
	input  [6:0]  iact_1_2_horiz_address_in_bits,
	output        iact_1_2_horiz_data_in_ready,
	input         iact_1_2_horiz_data_in_valid,         
	input  [11:0] iact_1_2_horiz_data_in_bits,          
	// dst port                                                    
	input         iact_1_2_PE_address_out_ready,        
	output        iact_1_2_PE_address_out_valid,         
	output [6:0]  iact_1_2_PE_address_out_bits,        
	input         iact_1_2_PE_data_out_ready,
	output        iact_1_2_PE_data_out_valid,
	output [11:0] iact_1_2_PE_data_out_bits,
						 
	input		  iact_1_2_north_address_out_ready,
	output        iact_1_2_north_address_out_valid,
	output [6:0]  iact_1_2_north_address_out_bits,
	input		  iact_1_2_north_data_out_ready,
	output        iact_1_2_north_data_out_valid,
	output [11:0] iact_1_2_north_data_out_bits,
						 
	input         iact_1_2_south_address_out_ready, 
	output        iact_1_2_south_address_out_valid,  
	output [6:0]  iact_1_2_south_address_out_bits, 
	input         iact_1_2_south_data_out_ready,
	output        iact_1_2_south_data_out_valid,
	output [11:0] iact_1_2_south_data_out_bits,
						 
	input         iact_1_2_horiz_address_out_ready, 
	output        iact_1_2_horiz_address_out_valid,  
	output [6:0]  iact_1_2_horiz_address_out_bits, 
	input         iact_1_2_horiz_data_out_ready,
	output        iact_1_2_horiz_data_out_valid,
	output [11:0] iact_1_2_horiz_data_out_bits,
	
	
	// ----------- iact router 2_0 ----------- //
	// src port
	output        iact_2_0_GLB_address_in_ready,
	input         iact_2_0_GLB_address_in_valid,
	input  [6:0]  iact_2_0_GLB_address_in_bits,
	output        iact_2_0_GLB_data_in_ready,
	input         iact_2_0_GLB_data_in_valid,
	input  [11:0] iact_2_0_GLB_data_in_bits,
						 
	output        iact_2_0_north_address_in_ready,
	input         iact_2_0_north_address_in_valid,
	input  [6:0]  iact_2_0_north_address_in_bits,
	output        iact_2_0_north_data_in_ready,
	input         iact_2_0_north_data_in_valid,
	input  [11:0] iact_2_0_north_data_in_bits,
						 
	output        iact_2_0_south_address_in_ready,
	input         iact_2_0_south_address_in_valid,
	input  [6:0]  iact_2_0_south_address_in_bits,
	output        iact_2_0_south_data_in_ready,
	input         iact_2_0_south_data_in_valid,
	input  [11:0] iact_2_0_south_data_in_bits,
						 
	output        iact_2_0_horiz_address_in_ready,
	input         iact_2_0_horiz_address_in_valid,
	input  [6:0]  iact_2_0_horiz_address_in_bits,
	output        iact_2_0_horiz_data_in_ready,
	input         iact_2_0_horiz_data_in_valid,         
	input  [11:0] iact_2_0_horiz_data_in_bits,          
	// dst port                                             
	input         iact_2_0_PE_address_out_ready,        
	output        iact_2_0_PE_address_out_valid,         
	output [6:0]  iact_2_0_PE_address_out_bits,        
	input         iact_2_0_PE_data_out_ready,
	output        iact_2_0_PE_data_out_valid,
	output [11:0] iact_2_0_PE_data_out_bits,
						 
	input		  iact_2_0_north_address_out_ready,
	output        iact_2_0_north_address_out_valid,
	output [6:0]  iact_2_0_north_address_out_bits,
	input		  iact_2_0_north_data_out_ready,
	output        iact_2_0_north_data_out_valid,
	output [11:0] iact_2_0_north_data_out_bits,
						 
	input         iact_2_0_south_address_out_ready, 
	output        iact_2_0_south_address_out_valid,  
	output [6:0]  iact_2_0_south_address_out_bits, 
	input         iact_2_0_south_data_out_ready,
	output        iact_2_0_south_data_out_valid,
	output [11:0] iact_2_0_south_data_out_bits,
						 
	input         iact_2_0_horiz_address_out_ready, 
	output        iact_2_0_horiz_address_out_valid,  
	output [6:0]  iact_2_0_horiz_address_out_bits, 
	input         iact_2_0_horiz_data_out_ready,
	output        iact_2_0_horiz_data_out_valid,
	output [11:0] iact_2_0_horiz_data_out_bits,
	
	
	// ----------- iact router 2_1 ----------- //
	// src port
	output        iact_2_1_GLB_address_in_ready,
	input         iact_2_1_GLB_address_in_valid,
	input  [6:0]  iact_2_1_GLB_address_in_bits,
	output        iact_2_1_GLB_data_in_ready,
	input         iact_2_1_GLB_data_in_valid,
	input  [11:0] iact_2_1_GLB_data_in_bits,
						 
	output        iact_2_1_north_address_in_ready,
	input         iact_2_1_north_address_in_valid,
	input  [6:0]  iact_2_1_north_address_in_bits,
	output        iact_2_1_north_data_in_ready,
	input         iact_2_1_north_data_in_valid,
	input  [11:0] iact_2_1_north_data_in_bits,
						 
	output        iact_2_1_south_address_in_ready,
	input         iact_2_1_south_address_in_valid,
	input  [6:0]  iact_2_1_south_address_in_bits,
	output        iact_2_1_south_data_in_ready,
	input         iact_2_1_south_data_in_valid,
	input  [11:0] iact_2_1_south_data_in_bits,
						 
	output        iact_2_1_horiz_address_in_ready,
	input         iact_2_1_horiz_address_in_valid,
	input  [6:0]  iact_2_1_horiz_address_in_bits,
	output        iact_2_1_horiz_data_in_ready,
	input         iact_2_1_horiz_data_in_valid,         
	input  [11:0] iact_2_1_horiz_data_in_bits,          
	// dst port                                           
	input         iact_2_1_PE_address_out_ready,        
	output        iact_2_1_PE_address_out_valid,         
	output [6:0]  iact_2_1_PE_address_out_bits,        
	input         iact_2_1_PE_data_out_ready,
	output        iact_2_1_PE_data_out_valid,
	output [11:0] iact_2_1_PE_data_out_bits,
						 
	input		  iact_2_1_north_address_out_ready,
	output        iact_2_1_north_address_out_valid,
	output [6:0]  iact_2_1_north_address_out_bits,
	input		  iact_2_1_north_data_out_ready,
	output        iact_2_1_north_data_out_valid,
	output [11:0] iact_2_1_north_data_out_bits,
						 
	input         iact_2_1_south_address_out_ready, 
	output        iact_2_1_south_address_out_valid,  
	output [6:0]  iact_2_1_south_address_out_bits, 
	input         iact_2_1_south_data_out_ready,
	output        iact_2_1_south_data_out_valid,
	output [11:0] iact_2_1_south_data_out_bits,
						 
	input         iact_2_1_horiz_address_out_ready, 
	output        iact_2_1_horiz_address_out_valid,  
	output [6:0]  iact_2_1_horiz_address_out_bits, 
	input         iact_2_1_horiz_data_out_ready,
	output        iact_2_1_horiz_data_out_valid,
	output [11:0] iact_2_1_horiz_data_out_bits,
	
	
	// ----------- iact router 2_2 ----------- //
	// src port
	output        iact_2_2_GLB_address_in_ready,
	input         iact_2_2_GLB_address_in_valid,
	input  [6:0]  iact_2_2_GLB_address_in_bits,
	output        iact_2_2_GLB_data_in_ready,
	input         iact_2_2_GLB_data_in_valid,
	input  [11:0] iact_2_2_GLB_data_in_bits,
						 
	output        iact_2_2_north_address_in_ready,
	input         iact_2_2_north_address_in_valid,
	input  [6:0]  iact_2_2_north_address_in_bits,
	output        iact_2_2_north_data_in_ready,
	input         iact_2_2_north_data_in_valid,
	input  [11:0] iact_2_2_north_data_in_bits,
						 
	output        iact_2_2_south_address_in_ready,
	input         iact_2_2_south_address_in_valid,
	input  [6:0]  iact_2_2_south_address_in_bits,
	output        iact_2_2_south_data_in_ready,
	input         iact_2_2_south_data_in_valid,
	input  [11:0] iact_2_2_south_data_in_bits,
						 
	output        iact_2_2_horiz_address_in_ready,
	input         iact_2_2_horiz_address_in_valid,
	input  [6:0]  iact_2_2_horiz_address_in_bits,
	output        iact_2_2_horiz_data_in_ready,
	input         iact_2_2_horiz_data_in_valid,         
	input  [11:0] iact_2_2_horiz_data_in_bits,          
	// dst port                                         
	input         iact_2_2_PE_address_out_ready,        
	output        iact_2_2_PE_address_out_valid,         
	output [6:0]  iact_2_2_PE_address_out_bits,        
	input         iact_2_2_PE_data_out_ready,
	output        iact_2_2_PE_data_out_valid,
	output [11:0] iact_2_2_PE_data_out_bits,
						 
	input		  iact_2_2_north_address_out_ready,
	output        iact_2_2_north_address_out_valid,
	output [6:0]  iact_2_2_north_address_out_bits,
	input		  iact_2_2_north_data_out_ready,
	output        iact_2_2_north_data_out_valid,
	output [11:0] iact_2_2_north_data_out_bits,
						 
	input         iact_2_2_south_address_out_ready, 
	output        iact_2_2_south_address_out_valid,  
	output [6:0]  iact_2_2_south_address_out_bits, 
	input         iact_2_2_south_data_out_ready,
	output        iact_2_2_south_data_out_valid,
	output [11:0] iact_2_2_south_data_out_bits,
						 
	input         iact_2_2_horiz_address_out_ready, 
	output        iact_2_2_horiz_address_out_valid,  
	output [6:0]  iact_2_2_horiz_address_out_bits, 
	input         iact_2_2_horiz_data_out_ready,
	output        iact_2_2_horiz_data_out_valid,
	output [11:0] iact_2_2_horiz_data_out_bits,
	
	
	// ----------- weight router 0 ----------- //
	// src port
	output        weight_0_GLB_address_in_ready,
	input         weight_0_GLB_address_in_valid,
	input  [7:0]  weight_0_GLB_address_in_bits,
	output        weight_0_GLB_data_in_ready,                                         
	input         weight_0_GLB_data_in_valid,                                         
	input  [12:0] weight_0_GLB_data_in_bits,                                          
	                                                                                  
	output        weight_0_horiz_address_in_ready,                                    
	input         weight_0_horiz_address_in_valid,                                    
	input  [7:0]  weight_0_horiz_address_in_bits,
	output        weight_0_horiz_data_in_ready,
	input         weight_0_horiz_data_in_valid,
	input  [12:0] weight_0_horiz_data_in_bits,
	// dst port     
	output        weight_0_PE_address_out_valid,
	output [7:0]  weight_0_PE_address_out_bits,
	output        weight_0_PE_data_out_valid,
	output [12:0] weight_0_PE_data_out_bits,
	
	input         weight_0_horiz_address_out_ready,  
	output        weight_0_horiz_address_out_valid,  
	output [7:0]  weight_0_horiz_address_out_bits,
	input         weight_0_horiz_data_out_ready,
	output        weight_0_horiz_data_out_valid,
	output [12:0] weight_0_horiz_data_out_bits,
	
	// ----------- weight router 1 ----------- //
	// src port
	output        weight_1_GLB_address_in_ready,
	input         weight_1_GLB_address_in_valid,
	input  [7:0]  weight_1_GLB_address_in_bits,
	output        weight_1_GLB_data_in_ready,        
	input         weight_1_GLB_data_in_valid,        
	input  [12:0] weight_1_GLB_data_in_bits,         
	                                               
	output        weight_1_horiz_address_in_ready,   
	input         weight_1_horiz_address_in_valid,   
	input  [7:0]  weight_1_horiz_address_in_bits,
	output        weight_1_horiz_data_in_ready,
	input         weight_1_horiz_data_in_valid,
	input  [12:0] weight_1_horiz_data_in_bits,
	// dst port               
	output        weight_1_PE_address_out_valid,
	output [7:0]  weight_1_PE_address_out_bits,
	output        weight_1_PE_data_out_valid,
	output [12:0] weight_1_PE_data_out_bits,
						 
	input         weight_1_horiz_address_out_ready,  
	output        weight_1_horiz_address_out_valid,  
	output [7:0]  weight_1_horiz_address_out_bits,
	input         weight_1_horiz_data_out_ready,
	output        weight_1_horiz_data_out_valid,
	output [12:0] weight_1_horiz_data_out_bits,
	
	// ----------- weight router 2 ----------- //
	// src port
	output        weight_2_GLB_address_in_ready,
	input         weight_2_GLB_address_in_valid,
	input  [7:0]  weight_2_GLB_address_in_bits,
	output        weight_2_GLB_data_in_ready,      
	input         weight_2_GLB_data_in_valid,      
	input  [12:0] weight_2_GLB_data_in_bits,       
	                                              
	output        weight_2_horiz_address_in_ready, 
	input         weight_2_horiz_address_in_valid, 
	input  [7:0]  weight_2_horiz_address_in_bits,
	output        weight_2_horiz_data_in_ready,
	input         weight_2_horiz_data_in_valid,
	input  [12:0] weight_2_horiz_data_in_bits,
	// dst port              
	output        weight_2_PE_address_out_valid,
	output [7:0]  weight_2_PE_address_out_bits,
	output        weight_2_PE_data_out_valid,
	output [12:0] weight_2_PE_data_out_bits,
						 
	input         weight_2_horiz_address_out_ready,
	output        weight_2_horiz_address_out_valid,
	output [7:0]  weight_2_horiz_address_out_bits,
	input         weight_2_horiz_data_out_ready,
	output        weight_2_horiz_data_out_valid,
	output [12:0] weight_2_horiz_data_out_bits,
	
	// ----------- psum router 0 ----------- //
	// src port
	output        		psum_0_PE_in_ready,
	input         		psum_0_PE_in_valid,
	input signed [20:0] psum_0_PE_in_bits,
	output        		psum_0_GLB_in_ready,
	input         		psum_0_GLB_in_valid,
	input signed [20:0] psum_0_GLB_in_bits,
	output        		psum_0_north_in_ready,
	input         		psum_0_north_in_valid,
	input signed [20:0] psum_0_north_in_bits,
	// dst port 
	input         		psum_0_PE_out_ready,
	output        		psum_0_PE_out_valid,
	output signed [20:0]psum_0_PE_out_bits,
	input         		psum_0_GLB_out_ready,
	output        		psum_0_GLB_out_valid,
	output signed [20:0]psum_0_GLB_out_bits,
	input        		psum_0_south_out_ready,
	output        		psum_0_south_out_valid,
	output signed [20:0]psum_0_south_out_bits,
	
	// ----------- psum router 1 ----------- //
	// src port
	output        		psum_1_PE_in_ready,
	input         		psum_1_PE_in_valid,
	input signed [20:0] psum_1_PE_in_bits,
	output        		psum_1_GLB_in_ready,
	input         		psum_1_GLB_in_valid,
	input signed [20:0] psum_1_GLB_in_bits,
	output        		psum_1_north_in_ready,
	input         		psum_1_north_in_valid,
	input signed [20:0] psum_1_north_in_bits,
	// dst port              
	input         		psum_1_PE_out_ready,
	output        		psum_1_PE_out_valid,
	output signed [20:0]psum_1_PE_out_bits,
	input         		psum_1_GLB_out_ready,
	output        		psum_1_GLB_out_valid,
	output signed [20:0]psum_1_GLB_out_bits,
	input        		psum_1_south_out_ready,
	output        		psum_1_south_out_valid,
	output signed [20:0]psum_1_south_out_bits,
	
	// ----------- psum router 2 ----------- //
	// src port
	output        		psum_2_PE_in_ready,
	input         		psum_2_PE_in_valid,
	input signed [20:0] psum_2_PE_in_bits,
	output        		psum_2_GLB_in_ready,
	input         		psum_2_GLB_in_valid,
	input signed [20:0] psum_2_GLB_in_bits,
	output        		psum_2_north_in_ready,
	input         		psum_2_north_in_valid,
	input signed [20:0] psum_2_north_in_bits,
	// dst port              
	input         		psum_2_PE_out_ready,
	output        		psum_2_PE_out_valid,
	output signed [20:0]psum_2_PE_out_bits,
	input         		psum_2_GLB_out_ready,
	output        		psum_2_GLB_out_valid,
	output signed [20:0]psum_2_GLB_out_bits,
	input        		psum_2_south_out_ready,
	output        		psum_2_south_out_valid,
	output signed [20:0]psum_2_south_out_bits
	
);

Iact_Router Iact_Router_0_0 ( 
	.GLB_address_in_ready   (iact_0_0_GLB_address_in_ready   	),
	.GLB_address_in_valid   (iact_0_0_GLB_address_in_valid   	),
	.GLB_address_in         (iact_0_0_GLB_address_in_bits		),
	.GLB_data_in_ready      (iact_0_0_GLB_data_in_ready      	),
	.GLB_data_in_valid      (iact_0_0_GLB_data_in_valid      	),
	.GLB_data_in	        (iact_0_0_GLB_data_in_bits			),
	.north_address_in_ready (iact_0_0_north_address_in_ready 	),
	.north_address_in_valid (iact_0_0_north_address_in_valid 	),
	.north_address_in       (iact_0_0_north_address_in_bits		),
	.north_data_in_ready    (iact_0_0_north_data_in_ready    	),
	.north_data_in_valid    (iact_0_0_north_data_in_valid    	),
	.north_data_in	        (iact_0_0_north_data_in_bits		),
	.south_address_in_ready (iact_0_0_south_address_in_ready 	),
	.south_address_in_valid (iact_0_0_south_address_in_valid 	),
	.south_address_in       (iact_0_0_south_address_in_bits		),
	.south_data_in_ready    (iact_0_0_south_data_in_ready    	),
	.south_data_in_valid    (iact_0_0_south_data_in_valid    	),
	.south_data_in	        (iact_0_0_south_data_in_bits		),
	.horiz_address_in_ready (iact_0_0_horiz_address_in_ready 	),
	.horiz_address_in_valid (iact_0_0_horiz_address_in_valid 	),
	.horiz_address_in       (iact_0_0_horiz_address_in_bits		),
	.horiz_data_in_ready    (iact_0_0_horiz_data_in_ready    	),
	.horiz_data_in_valid    (iact_0_0_horiz_data_in_valid    	),
	.horiz_data_in          (iact_0_0_horiz_data_in_bits	  	),
	.PE_address_out_ready   (iact_0_0_PE_address_out_ready   	),
	.PE_address_out_valid   (iact_0_0_PE_address_out_valid   	),
	.PE_address_out         (iact_0_0_PE_address_out_bits	    ),
	.PE_data_out_ready      (iact_0_0_PE_data_out_ready      	),
	.PE_data_out_valid      (iact_0_0_PE_data_out_valid      	),
	.PE_data_out            (iact_0_0_PE_data_out_bits	    	),
	.north_address_out_ready(iact_0_0_north_address_out_ready	),
	.north_address_out_valid(iact_0_0_north_address_out_valid	),
	.north_address_out      (iact_0_0_north_address_out_bits	),
	.north_data_out_ready	(iact_0_0_north_data_out_ready		),
	.north_data_out_valid   (iact_0_0_north_data_out_valid   	),
	.north_data_out         (iact_0_0_north_data_out_bits	    ),
	.south_address_out_ready(iact_0_0_south_address_out_ready	),
	.south_address_out_valid(iact_0_0_south_address_out_valid	),
	.south_address_out      (iact_0_0_south_address_out_bits	),
	.south_data_out_ready   (iact_0_0_south_data_out_ready   	),
	.south_data_out_valid   (iact_0_0_south_data_out_valid   	),
	.south_data_out         (iact_0_0_south_data_out_bits	    ),
	.horiz_address_out_ready(iact_0_0_horiz_address_out_ready	),
	.horiz_address_out_valid(iact_0_0_horiz_address_out_valid	),
	.horiz_address_out      (iact_0_0_horiz_address_out_bits	),
	.horiz_data_out_ready   (iact_0_0_horiz_data_out_ready   	),
	.horiz_data_out_valid   (iact_0_0_horiz_data_out_valid   	),
	.horiz_data_out         (iact_0_0_horiz_data_out_bits	    ),
	.data_in_sel            (iact_0_data_in_sel            		),
	.data_out_sel			(iact_0_data_out_sel				)
);

Iact_Router Iact_Router_0_1 ( 
	.GLB_address_in_ready   (iact_0_1_GLB_address_in_ready   	),
	.GLB_address_in_valid   (iact_0_1_GLB_address_in_valid   	),
	.GLB_address_in         (iact_0_1_GLB_address_in_bits		),
	.GLB_data_in_ready      (iact_0_1_GLB_data_in_ready      	),
	.GLB_data_in_valid      (iact_0_1_GLB_data_in_valid      	),
	.GLB_data_in	        (iact_0_1_GLB_data_in_bits			),
	.north_address_in_ready (iact_0_1_north_address_in_ready 	),
	.north_address_in_valid (iact_0_1_north_address_in_valid 	),
	.north_address_in       (iact_0_1_north_address_in_bits		),
	.north_data_in_ready    (iact_0_1_north_data_in_ready    	),
	.north_data_in_valid    (iact_0_1_north_data_in_valid    	),
	.north_data_in	        (iact_0_1_north_data_in_bits		),
	.south_address_in_ready (iact_0_1_south_address_in_ready 	),
	.south_address_in_valid (iact_0_1_south_address_in_valid 	),
	.south_address_in       (iact_0_1_south_address_in_bits		),
	.south_data_in_ready    (iact_0_1_south_data_in_ready    	),
	.south_data_in_valid    (iact_0_1_south_data_in_valid    	),
	.south_data_in	        (iact_0_1_south_data_in_bits		),
	.horiz_address_in_ready (iact_0_1_horiz_address_in_ready 	),
	.horiz_address_in_valid (iact_0_1_horiz_address_in_valid 	),
	.horiz_address_in       (iact_0_1_horiz_address_in_bits		),
	.horiz_data_in_ready    (iact_0_1_horiz_data_in_ready    	),
	.horiz_data_in_valid    (iact_0_1_horiz_data_in_valid    	),
	.horiz_data_in          (iact_0_1_horiz_data_in_bits	  	),
	.PE_address_out_ready   (iact_0_1_PE_address_out_ready   	),
	.PE_address_out_valid   (iact_0_1_PE_address_out_valid   	),
	.PE_address_out         (iact_0_1_PE_address_out_bits	    ),
	.PE_data_out_ready      (iact_0_1_PE_data_out_ready      	),
	.PE_data_out_valid      (iact_0_1_PE_data_out_valid      	),
	.PE_data_out            (iact_0_1_PE_data_out_bits	    	),
	.north_address_out_ready(iact_0_1_north_address_out_ready	),
	.north_address_out_valid(iact_0_1_north_address_out_valid	),
	.north_address_out      (iact_0_1_north_address_out_bits	),
	.north_data_out_ready	(iact_0_1_north_data_out_ready		),
	.north_data_out_valid   (iact_0_1_north_data_out_valid   	),
	.north_data_out         (iact_0_1_north_data_out_bits	    ),
	.south_address_out_ready(iact_0_1_south_address_out_ready	),
	.south_address_out_valid(iact_0_1_south_address_out_valid	),
	.south_address_out      (iact_0_1_south_address_out_bits	),
	.south_data_out_ready   (iact_0_1_south_data_out_ready   	),
	.south_data_out_valid   (iact_0_1_south_data_out_valid   	),
	.south_data_out         (iact_0_1_south_data_out_bits	    ),
	.horiz_address_out_ready(iact_0_1_horiz_address_out_ready	),
	.horiz_address_out_valid(iact_0_1_horiz_address_out_valid	),
	.horiz_address_out      (iact_0_1_horiz_address_out_bits	),
	.horiz_data_out_ready   (iact_0_1_horiz_data_out_ready   	),
	.horiz_data_out_valid   (iact_0_1_horiz_data_out_valid   	),
	.horiz_data_out         (iact_0_1_horiz_data_out_bits	    ),
	.data_in_sel            (iact_0_data_in_sel            		),
	.data_out_sel			(iact_0_data_out_sel				)
);

Iact_Router Iact_Router_0_2 ( 
	.GLB_address_in_ready   (iact_0_2_GLB_address_in_ready   	),
	.GLB_address_in_valid   (iact_0_2_GLB_address_in_valid   	),
	.GLB_address_in         (iact_0_2_GLB_address_in_bits		),
	.GLB_data_in_ready      (iact_0_2_GLB_data_in_ready      	),
	.GLB_data_in_valid      (iact_0_2_GLB_data_in_valid      	),
	.GLB_data_in	        (iact_0_2_GLB_data_in_bits			),
	.north_address_in_ready (iact_0_2_north_address_in_ready 	),
	.north_address_in_valid (iact_0_2_north_address_in_valid 	),
	.north_address_in       (iact_0_2_north_address_in_bits		),
	.north_data_in_ready    (iact_0_2_north_data_in_ready    	),
	.north_data_in_valid    (iact_0_2_north_data_in_valid    	),
	.north_data_in	        (iact_0_2_north_data_in_bits		),
	.south_address_in_ready (iact_0_2_south_address_in_ready 	),
	.south_address_in_valid (iact_0_2_south_address_in_valid 	),
	.south_address_in       (iact_0_2_south_address_in_bits		),
	.south_data_in_ready    (iact_0_2_south_data_in_ready    	),
	.south_data_in_valid    (iact_0_2_south_data_in_valid    	),
	.south_data_in	        (iact_0_2_south_data_in_bits		),
	.horiz_address_in_ready (iact_0_2_horiz_address_in_ready 	),
	.horiz_address_in_valid (iact_0_2_horiz_address_in_valid 	),
	.horiz_address_in       (iact_0_2_horiz_address_in_bits		),
	.horiz_data_in_ready    (iact_0_2_horiz_data_in_ready    	),
	.horiz_data_in_valid    (iact_0_2_horiz_data_in_valid    	),
	.horiz_data_in          (iact_0_2_horiz_data_in_bits	  	),
	.PE_address_out_ready   (iact_0_2_PE_address_out_ready   	),
	.PE_address_out_valid   (iact_0_2_PE_address_out_valid   	),
	.PE_address_out         (iact_0_2_PE_address_out_bits	    ),
	.PE_data_out_ready      (iact_0_2_PE_data_out_ready      	),
	.PE_data_out_valid      (iact_0_2_PE_data_out_valid      	),
	.PE_data_out            (iact_0_2_PE_data_out_bits	    	),
	.north_address_out_ready(iact_0_2_north_address_out_ready	),
	.north_address_out_valid(iact_0_2_north_address_out_valid	),
	.north_address_out      (iact_0_2_north_address_out_bits	),
	.north_data_out_ready	(iact_0_2_north_data_out_ready		),
	.north_data_out_valid   (iact_0_2_north_data_out_valid   	),
	.north_data_out         (iact_0_2_north_data_out_bits	    ),
	.south_address_out_ready(iact_0_2_south_address_out_ready	),
	.south_address_out_valid(iact_0_2_south_address_out_valid	),
	.south_address_out      (iact_0_2_south_address_out_bits	),
	.south_data_out_ready   (iact_0_2_south_data_out_ready   	),
	.south_data_out_valid   (iact_0_2_south_data_out_valid   	),
	.south_data_out         (iact_0_2_south_data_out_bits	    ),
	.horiz_address_out_ready(iact_0_2_horiz_address_out_ready	),
	.horiz_address_out_valid(iact_0_2_horiz_address_out_valid	),
	.horiz_address_out      (iact_0_2_horiz_address_out_bits	),
	.horiz_data_out_ready   (iact_0_2_horiz_data_out_ready   	),
	.horiz_data_out_valid   (iact_0_2_horiz_data_out_valid   	),
	.horiz_data_out         (iact_0_2_horiz_data_out_bits	    ),
	.data_in_sel            (iact_0_data_in_sel            		),
	.data_out_sel			(iact_0_data_out_sel				)
);


Iact_Router Iact_Router_1_0 ( 
	.GLB_address_in_ready   (iact_1_0_GLB_address_in_ready   	),
	.GLB_address_in_valid   (iact_1_0_GLB_address_in_valid   	),
	.GLB_address_in         (iact_1_0_GLB_address_in_bits		),
	.GLB_data_in_ready      (iact_1_0_GLB_data_in_ready      	),
	.GLB_data_in_valid      (iact_1_0_GLB_data_in_valid      	),
	.GLB_data_in	        (iact_1_0_GLB_data_in_bits			),
	.north_address_in_ready (iact_1_0_north_address_in_ready 	),
	.north_address_in_valid (iact_1_0_north_address_in_valid 	),
	.north_address_in       (iact_1_0_north_address_in_bits		),
	.north_data_in_ready    (iact_1_0_north_data_in_ready    	),
	.north_data_in_valid    (iact_1_0_north_data_in_valid    	),
	.north_data_in	        (iact_1_0_north_data_in_bits		),
	.south_address_in_ready (iact_1_0_south_address_in_ready 	),
	.south_address_in_valid (iact_1_0_south_address_in_valid 	),
	.south_address_in       (iact_1_0_south_address_in_bits		),
	.south_data_in_ready    (iact_1_0_south_data_in_ready    	),
	.south_data_in_valid    (iact_1_0_south_data_in_valid    	),
	.south_data_in	        (iact_1_0_south_data_in_bits		),
	.horiz_address_in_ready (iact_1_0_horiz_address_in_ready 	),
	.horiz_address_in_valid (iact_1_0_horiz_address_in_valid 	),
	.horiz_address_in       (iact_1_0_horiz_address_in_bits		),
	.horiz_data_in_ready    (iact_1_0_horiz_data_in_ready    	),
	.horiz_data_in_valid    (iact_1_0_horiz_data_in_valid    	),
	.horiz_data_in          (iact_1_0_horiz_data_in_bits	  	),
	.PE_address_out_ready   (iact_1_0_PE_address_out_ready   	),
	.PE_address_out_valid   (iact_1_0_PE_address_out_valid   	),
	.PE_address_out         (iact_1_0_PE_address_out_bits	    ),
	.PE_data_out_ready      (iact_1_0_PE_data_out_ready      	),
	.PE_data_out_valid      (iact_1_0_PE_data_out_valid      	),
	.PE_data_out            (iact_1_0_PE_data_out_bits	    	),
	.north_address_out_ready(iact_1_0_north_address_out_ready	),
	.north_address_out_valid(iact_1_0_north_address_out_valid	),
	.north_address_out      (iact_1_0_north_address_out_bits	),
	.north_data_out_ready	(iact_1_0_north_data_out_ready		),
	.north_data_out_valid   (iact_1_0_north_data_out_valid   	),
	.north_data_out         (iact_1_0_north_data_out_bits	    ),
	.south_address_out_ready(iact_1_0_south_address_out_ready	),
	.south_address_out_valid(iact_1_0_south_address_out_valid	),
	.south_address_out      (iact_1_0_south_address_out_bits	),
	.south_data_out_ready   (iact_1_0_south_data_out_ready   	),
	.south_data_out_valid   (iact_1_0_south_data_out_valid   	),
	.south_data_out         (iact_1_0_south_data_out_bits	    ),
	.horiz_address_out_ready(iact_1_0_horiz_address_out_ready	),
	.horiz_address_out_valid(iact_1_0_horiz_address_out_valid	),
	.horiz_address_out      (iact_1_0_horiz_address_out_bits	),
	.horiz_data_out_ready   (iact_1_0_horiz_data_out_ready   	),
	.horiz_data_out_valid   (iact_1_0_horiz_data_out_valid   	),
	.horiz_data_out         (iact_1_0_horiz_data_out_bits	    ),
	.data_in_sel            (iact_1_data_in_sel            		),
	.data_out_sel			(iact_1_data_out_sel				)
);


Iact_Router Iact_Router_1_1 ( 
	.GLB_address_in_ready   (iact_1_1_GLB_address_in_ready   	),
	.GLB_address_in_valid   (iact_1_1_GLB_address_in_valid   	),
	.GLB_address_in         (iact_1_1_GLB_address_in_bits		),
	.GLB_data_in_ready      (iact_1_1_GLB_data_in_ready      	),
	.GLB_data_in_valid      (iact_1_1_GLB_data_in_valid      	),
	.GLB_data_in	        (iact_1_1_GLB_data_in_bits			),
	.north_address_in_ready (iact_1_1_north_address_in_ready 	),
	.north_address_in_valid (iact_1_1_north_address_in_valid 	),
	.north_address_in       (iact_1_1_north_address_in_bits		),
	.north_data_in_ready    (iact_1_1_north_data_in_ready    	),
	.north_data_in_valid    (iact_1_1_north_data_in_valid    	),
	.north_data_in	        (iact_1_1_north_data_in_bits		),
	.south_address_in_ready (iact_1_1_south_address_in_ready 	),
	.south_address_in_valid (iact_1_1_south_address_in_valid 	),
	.south_address_in       (iact_1_1_south_address_in_bits		),
	.south_data_in_ready    (iact_1_1_south_data_in_ready    	),
	.south_data_in_valid    (iact_1_1_south_data_in_valid    	),
	.south_data_in	        (iact_1_1_south_data_in_bits		),
	.horiz_address_in_ready (iact_1_1_horiz_address_in_ready 	),
	.horiz_address_in_valid (iact_1_1_horiz_address_in_valid 	),
	.horiz_address_in       (iact_1_1_horiz_address_in_bits		),
	.horiz_data_in_ready    (iact_1_1_horiz_data_in_ready    	),
	.horiz_data_in_valid    (iact_1_1_horiz_data_in_valid    	),
	.horiz_data_in          (iact_1_1_horiz_data_in_bits	  	),
	.PE_address_out_ready   (iact_1_1_PE_address_out_ready   	),
	.PE_address_out_valid   (iact_1_1_PE_address_out_valid   	),
	.PE_address_out         (iact_1_1_PE_address_out_bits	    ),
	.PE_data_out_ready      (iact_1_1_PE_data_out_ready      	),
	.PE_data_out_valid      (iact_1_1_PE_data_out_valid      	),
	.PE_data_out            (iact_1_1_PE_data_out_bits	    	),
	.north_address_out_ready(iact_1_1_north_address_out_ready	),
	.north_address_out_valid(iact_1_1_north_address_out_valid	),
	.north_address_out      (iact_1_1_north_address_out_bits	),
	.north_data_out_ready	(iact_1_1_north_data_out_ready		),
	.north_data_out_valid   (iact_1_1_north_data_out_valid   	),
	.north_data_out         (iact_1_1_north_data_out_bits	    ),
	.south_address_out_ready(iact_1_1_south_address_out_ready	),
	.south_address_out_valid(iact_1_1_south_address_out_valid	),
	.south_address_out      (iact_1_1_south_address_out_bits	),
	.south_data_out_ready   (iact_1_1_south_data_out_ready   	),
	.south_data_out_valid   (iact_1_1_south_data_out_valid   	),
	.south_data_out         (iact_1_1_south_data_out_bits	    ),
	.horiz_address_out_ready(iact_1_1_horiz_address_out_ready	),
	.horiz_address_out_valid(iact_1_1_horiz_address_out_valid	),
	.horiz_address_out      (iact_1_1_horiz_address_out_bits	),
	.horiz_data_out_ready   (iact_1_1_horiz_data_out_ready   	),
	.horiz_data_out_valid   (iact_1_1_horiz_data_out_valid   	),
	.horiz_data_out         (iact_1_1_horiz_data_out_bits	    ),
	.data_in_sel            (iact_1_data_in_sel            		),
	.data_out_sel			(iact_1_data_out_sel				)
);


Iact_Router Iact_Router_1_2 ( 
	.GLB_address_in_ready   (iact_1_2_GLB_address_in_ready   	),
	.GLB_address_in_valid   (iact_1_2_GLB_address_in_valid   	),
	.GLB_address_in         (iact_1_2_GLB_address_in_bits		),
	.GLB_data_in_ready      (iact_1_2_GLB_data_in_ready      	),
	.GLB_data_in_valid      (iact_1_2_GLB_data_in_valid      	),
	.GLB_data_in	        (iact_1_2_GLB_data_in_bits			),
	.north_address_in_ready (iact_1_2_north_address_in_ready 	),
	.north_address_in_valid (iact_1_2_north_address_in_valid 	),
	.north_address_in       (iact_1_2_north_address_in_bits		),
	.north_data_in_ready    (iact_1_2_north_data_in_ready    	),
	.north_data_in_valid    (iact_1_2_north_data_in_valid    	),
	.north_data_in	        (iact_1_2_north_data_in_bits		),
	.south_address_in_ready (iact_1_2_south_address_in_ready 	),
	.south_address_in_valid (iact_1_2_south_address_in_valid 	),
	.south_address_in       (iact_1_2_south_address_in_bits		),
	.south_data_in_ready    (iact_1_2_south_data_in_ready    	),
	.south_data_in_valid    (iact_1_2_south_data_in_valid    	),
	.south_data_in	        (iact_1_2_south_data_in_bits		),
	.horiz_address_in_ready (iact_1_2_horiz_address_in_ready 	),
	.horiz_address_in_valid (iact_1_2_horiz_address_in_valid 	),
	.horiz_address_in       (iact_1_2_horiz_address_in_bits		),
	.horiz_data_in_ready    (iact_1_2_horiz_data_in_ready    	),
	.horiz_data_in_valid    (iact_1_2_horiz_data_in_valid    	),
	.horiz_data_in          (iact_1_2_horiz_data_in_bits	  	),
	.PE_address_out_ready   (iact_1_2_PE_address_out_ready   	),
	.PE_address_out_valid   (iact_1_2_PE_address_out_valid   	),
	.PE_address_out         (iact_1_2_PE_address_out_bits	    ),
	.PE_data_out_ready      (iact_1_2_PE_data_out_ready      	),
	.PE_data_out_valid      (iact_1_2_PE_data_out_valid      	),
	.PE_data_out            (iact_1_2_PE_data_out_bits	    	),
	.north_address_out_ready(iact_1_2_north_address_out_ready	),
	.north_address_out_valid(iact_1_2_north_address_out_valid	),
	.north_address_out      (iact_1_2_north_address_out_bits	),
	.north_data_out_ready	(iact_1_2_north_data_out_ready		),
	.north_data_out_valid   (iact_1_2_north_data_out_valid   	),
	.north_data_out         (iact_1_2_north_data_out_bits	    ),
	.south_address_out_ready(iact_1_2_south_address_out_ready	),
	.south_address_out_valid(iact_1_2_south_address_out_valid	),
	.south_address_out      (iact_1_2_south_address_out_bits	),
	.south_data_out_ready   (iact_1_2_south_data_out_ready   	),
	.south_data_out_valid   (iact_1_2_south_data_out_valid   	),
	.south_data_out         (iact_1_2_south_data_out_bits	    ),
	.horiz_address_out_ready(iact_1_2_horiz_address_out_ready	),
	.horiz_address_out_valid(iact_1_2_horiz_address_out_valid	),
	.horiz_address_out      (iact_1_2_horiz_address_out_bits	),
	.horiz_data_out_ready   (iact_1_2_horiz_data_out_ready   	),
	.horiz_data_out_valid   (iact_1_2_horiz_data_out_valid   	),
	.horiz_data_out         (iact_1_2_horiz_data_out_bits	    ),
	.data_in_sel            (iact_1_data_in_sel            		),
	.data_out_sel			(iact_1_data_out_sel				)
);


Iact_Router Iact_Router_2_0 ( 
	.GLB_address_in_ready   (iact_2_0_GLB_address_in_ready   	),
	.GLB_address_in_valid   (iact_2_0_GLB_address_in_valid   	),
	.GLB_address_in         (iact_2_0_GLB_address_in_bits		),
	.GLB_data_in_ready      (iact_2_0_GLB_data_in_ready      	),
	.GLB_data_in_valid      (iact_2_0_GLB_data_in_valid      	),
	.GLB_data_in	        (iact_2_0_GLB_data_in_bits			),
	.north_address_in_ready (iact_2_0_north_address_in_ready 	),
	.north_address_in_valid (iact_2_0_north_address_in_valid 	),
	.north_address_in       (iact_2_0_north_address_in_bits		),
	.north_data_in_ready    (iact_2_0_north_data_in_ready    	),
	.north_data_in_valid    (iact_2_0_north_data_in_valid    	),
	.north_data_in	        (iact_2_0_north_data_in_bits		),
	.south_address_in_ready (iact_2_0_south_address_in_ready 	),
	.south_address_in_valid (iact_2_0_south_address_in_valid 	),
	.south_address_in       (iact_2_0_south_address_in_bits		),
	.south_data_in_ready    (iact_2_0_south_data_in_ready    	),
	.south_data_in_valid    (iact_2_0_south_data_in_valid    	),
	.south_data_in	        (iact_2_0_south_data_in_bits		),
	.horiz_address_in_ready (iact_2_0_horiz_address_in_ready 	),
	.horiz_address_in_valid (iact_2_0_horiz_address_in_valid 	),
	.horiz_address_in       (iact_2_0_horiz_address_in_bits		),
	.horiz_data_in_ready    (iact_2_0_horiz_data_in_ready    	),
	.horiz_data_in_valid    (iact_2_0_horiz_data_in_valid    	),
	.horiz_data_in          (iact_2_0_horiz_data_in_bits	  	),
	.PE_address_out_ready   (iact_2_0_PE_address_out_ready   	),
	.PE_address_out_valid   (iact_2_0_PE_address_out_valid   	),
	.PE_address_out         (iact_2_0_PE_address_out_bits	    ),
	.PE_data_out_ready      (iact_2_0_PE_data_out_ready      	),
	.PE_data_out_valid      (iact_2_0_PE_data_out_valid      	),
	.PE_data_out            (iact_2_0_PE_data_out_bits	    	),
	.north_address_out_ready(iact_2_0_north_address_out_ready	),
	.north_address_out_valid(iact_2_0_north_address_out_valid	),
	.north_address_out      (iact_2_0_north_address_out_bits	),
	.north_data_out_ready	(iact_2_0_north_data_out_ready		),
	.north_data_out_valid   (iact_2_0_north_data_out_valid   	),
	.north_data_out         (iact_2_0_north_data_out_bits	    ),
	.south_address_out_ready(iact_2_0_south_address_out_ready	),
	.south_address_out_valid(iact_2_0_south_address_out_valid	),
	.south_address_out      (iact_2_0_south_address_out_bits	),
	.south_data_out_ready   (iact_2_0_south_data_out_ready   	),
	.south_data_out_valid   (iact_2_0_south_data_out_valid   	),
	.south_data_out         (iact_2_0_south_data_out_bits	    ),
	.horiz_address_out_ready(iact_2_0_horiz_address_out_ready	),
	.horiz_address_out_valid(iact_2_0_horiz_address_out_valid	),
	.horiz_address_out      (iact_2_0_horiz_address_out_bits	),
	.horiz_data_out_ready   (iact_2_0_horiz_data_out_ready   	),
	.horiz_data_out_valid   (iact_2_0_horiz_data_out_valid   	),
	.horiz_data_out         (iact_2_0_horiz_data_out_bits	    ),
	.data_in_sel            (iact_2_data_in_sel           	 	),
	.data_out_sel			(iact_2_data_out_sel				)
);


Iact_Router Iact_Router_2_1 ( 
	.GLB_address_in_ready   (iact_2_1_GLB_address_in_ready   	),
	.GLB_address_in_valid   (iact_2_1_GLB_address_in_valid   	),
	.GLB_address_in         (iact_2_1_GLB_address_in_bits		),
	.GLB_data_in_ready      (iact_2_1_GLB_data_in_ready      	),
	.GLB_data_in_valid      (iact_2_1_GLB_data_in_valid      	),
	.GLB_data_in	        (iact_2_1_GLB_data_in_bits			),
	.north_address_in_ready (iact_2_1_north_address_in_ready 	),
	.north_address_in_valid (iact_2_1_north_address_in_valid 	),
	.north_address_in       (iact_2_1_north_address_in_bits		),
	.north_data_in_ready    (iact_2_1_north_data_in_ready    	),
	.north_data_in_valid    (iact_2_1_north_data_in_valid    	),
	.north_data_in	        (iact_2_1_north_data_in_bits		),
	.south_address_in_ready (iact_2_1_south_address_in_ready 	),
	.south_address_in_valid (iact_2_1_south_address_in_valid 	),
	.south_address_in       (iact_2_1_south_address_in_bits		),
	.south_data_in_ready    (iact_2_1_south_data_in_ready    	),
	.south_data_in_valid    (iact_2_1_south_data_in_valid    	),
	.south_data_in	        (iact_2_1_south_data_in_bits		),
	.horiz_address_in_ready (iact_2_1_horiz_address_in_ready 	),
	.horiz_address_in_valid (iact_2_1_horiz_address_in_valid 	),
	.horiz_address_in       (iact_2_1_horiz_address_in_bits		),
	.horiz_data_in_ready    (iact_2_1_horiz_data_in_ready    	),
	.horiz_data_in_valid    (iact_2_1_horiz_data_in_valid    	),
	.horiz_data_in          (iact_2_1_horiz_data_in_bits	  	),
	.PE_address_out_ready   (iact_2_1_PE_address_out_ready   	),
	.PE_address_out_valid   (iact_2_1_PE_address_out_valid   	),
	.PE_address_out         (iact_2_1_PE_address_out_bits	    ),
	.PE_data_out_ready      (iact_2_1_PE_data_out_ready      	),
	.PE_data_out_valid      (iact_2_1_PE_data_out_valid      	),
	.PE_data_out            (iact_2_1_PE_data_out_bits	    	),
	.north_address_out_ready(iact_2_1_north_address_out_ready	),
	.north_address_out_valid(iact_2_1_north_address_out_valid	),
	.north_address_out      (iact_2_1_north_address_out_bits	),
	.north_data_out_ready	(iact_2_1_north_data_out_ready		),
	.north_data_out_valid   (iact_2_1_north_data_out_valid   	),
	.north_data_out         (iact_2_1_north_data_out_bits	    ),
	.south_address_out_ready(iact_2_1_south_address_out_ready	),
	.south_address_out_valid(iact_2_1_south_address_out_valid	),
	.south_address_out      (iact_2_1_south_address_out_bits	),
	.south_data_out_ready   (iact_2_1_south_data_out_ready   	),
	.south_data_out_valid   (iact_2_1_south_data_out_valid   	),
	.south_data_out         (iact_2_1_south_data_out_bits	    ),
	.horiz_address_out_ready(iact_2_1_horiz_address_out_ready	),
	.horiz_address_out_valid(iact_2_1_horiz_address_out_valid	),
	.horiz_address_out      (iact_2_1_horiz_address_out_bits	),
	.horiz_data_out_ready   (iact_2_1_horiz_data_out_ready   	),
	.horiz_data_out_valid   (iact_2_1_horiz_data_out_valid   	),
	.horiz_data_out         (iact_2_1_horiz_data_out_bits	    ),
	.data_in_sel            (iact_2_data_in_sel            		),
	.data_out_sel			(iact_2_data_out_sel				)
);


Iact_Router Iact_Router_2_2 ( 
	.GLB_address_in_ready   (iact_2_2_GLB_address_in_ready   	),
	.GLB_address_in_valid   (iact_2_2_GLB_address_in_valid   	),
	.GLB_address_in         (iact_2_2_GLB_address_in_bits		),
	.GLB_data_in_ready      (iact_2_2_GLB_data_in_ready      	),
	.GLB_data_in_valid      (iact_2_2_GLB_data_in_valid      	),
	.GLB_data_in	        (iact_2_2_GLB_data_in_bits			),
	.north_address_in_ready (iact_2_2_north_address_in_ready 	),
	.north_address_in_valid (iact_2_2_north_address_in_valid 	),
	.north_address_in       (iact_2_2_north_address_in_bits		),
	.north_data_in_ready    (iact_2_2_north_data_in_ready    	),
	.north_data_in_valid    (iact_2_2_north_data_in_valid    	),
	.north_data_in	        (iact_2_2_north_data_in_bits		),
	.south_address_in_ready (iact_2_2_south_address_in_ready 	),
	.south_address_in_valid (iact_2_2_south_address_in_valid 	),
	.south_address_in       (iact_2_2_south_address_in_bits		),
	.south_data_in_ready    (iact_2_2_south_data_in_ready    	),
	.south_data_in_valid    (iact_2_2_south_data_in_valid    	),
	.south_data_in	        (iact_2_2_south_data_in_bits		),
	.horiz_address_in_ready (iact_2_2_horiz_address_in_ready 	),
	.horiz_address_in_valid (iact_2_2_horiz_address_in_valid 	),
	.horiz_address_in       (iact_2_2_horiz_address_in_bits		),
	.horiz_data_in_ready    (iact_2_2_horiz_data_in_ready    	),
	.horiz_data_in_valid    (iact_2_2_horiz_data_in_valid    	),
	.horiz_data_in          (iact_2_2_horiz_data_in_bits	  	),
	.PE_address_out_ready   (iact_2_2_PE_address_out_ready   	),
	.PE_address_out_valid   (iact_2_2_PE_address_out_valid   	),
	.PE_address_out         (iact_2_2_PE_address_out_bits	    ),
	.PE_data_out_ready      (iact_2_2_PE_data_out_ready      	),
	.PE_data_out_valid      (iact_2_2_PE_data_out_valid      	),
	.PE_data_out            (iact_2_2_PE_data_out_bits	    	),
	.north_address_out_ready(iact_2_2_north_address_out_ready	),
	.north_address_out_valid(iact_2_2_north_address_out_valid	),
	.north_address_out      (iact_2_2_north_address_out_bits	),
	.north_data_out_ready	(iact_2_2_north_data_out_ready		),
	.north_data_out_valid   (iact_2_2_north_data_out_valid   	),
	.north_data_out         (iact_2_2_north_data_out_bits	    ),
	.south_address_out_ready(iact_2_2_south_address_out_ready	),
	.south_address_out_valid(iact_2_2_south_address_out_valid	),
	.south_address_out      (iact_2_2_south_address_out_bits	),
	.south_data_out_ready   (iact_2_2_south_data_out_ready   	),
	.south_data_out_valid   (iact_2_2_south_data_out_valid   	),
	.south_data_out         (iact_2_2_south_data_out_bits	    ),
	.horiz_address_out_ready(iact_2_2_horiz_address_out_ready	),
	.horiz_address_out_valid(iact_2_2_horiz_address_out_valid	),
	.horiz_address_out      (iact_2_2_horiz_address_out_bits	),
	.horiz_data_out_ready   (iact_2_2_horiz_data_out_ready   	),
	.horiz_data_out_valid   (iact_2_2_horiz_data_out_valid   	),
	.horiz_data_out         (iact_2_2_horiz_data_out_bits	    ),
	.data_in_sel            (iact_2_data_in_sel            		),
	.data_out_sel			(iact_2_data_out_sel				)
);


Weight_Router Weight_Router_0 ( 
	.GLB_address_in_ready	(weight_0_GLB_address_in_ready	 	),
	.GLB_address_in_valid   (weight_0_GLB_address_in_valid   	),
	.GLB_address_in         (weight_0_GLB_address_in_bits		),
	.GLB_data_in_ready      (weight_0_GLB_data_in_ready      	),
	.GLB_data_in_valid      (weight_0_GLB_data_in_valid      	),
	.GLB_data_in            (weight_0_GLB_data_in_bits			),
	.horiz_address_in_ready (weight_0_horiz_address_in_ready 	),
	.horiz_address_in_valid (weight_0_horiz_address_in_valid 	),
	.horiz_address_in       (weight_0_horiz_address_in_bits		),
	.horiz_data_in_ready    (weight_0_horiz_data_in_ready    	),
	.horiz_data_in_valid    (weight_0_horiz_data_in_valid    	),
	.horiz_data_in          (weight_0_horiz_data_in_bits		),
	.PE_address_out_valid   (weight_0_PE_address_out_valid   	),
	.PE_address_out         (weight_0_PE_address_out_bits		),
	.PE_data_out_valid      (weight_0_PE_data_out_valid      	),
	.PE_data_out            (weight_0_PE_data_out_bits			),
	.horiz_address_out_ready(weight_0_horiz_address_out_ready	),
	.horiz_address_out_valid(weight_0_horiz_address_out_valid	),
	.horiz_address_out      (weight_0_horiz_address_out_bits	),
	.horiz_data_out_ready   (weight_0_horiz_data_out_ready   	),
	.horiz_data_out_valid   (weight_0_horiz_data_out_valid   	),
	.horiz_data_out         (weight_0_horiz_data_out_bits		),
	.data_in_sel            (weight_0_data_in_sel            	),
	.data_out_sel           (weight_0_data_out_sel           	)
);

Weight_Router Weight_Router_1 ( 
	.GLB_address_in_ready	(weight_1_GLB_address_in_ready	 	),
	.GLB_address_in_valid   (weight_1_GLB_address_in_valid   	),
	.GLB_address_in         (weight_1_GLB_address_in_bits		),
	.GLB_data_in_ready      (weight_1_GLB_data_in_ready      	),
	.GLB_data_in_valid      (weight_1_GLB_data_in_valid      	),
	.GLB_data_in            (weight_1_GLB_data_in_bits			),
	.horiz_address_in_ready (weight_1_horiz_address_in_ready 	),
	.horiz_address_in_valid (weight_1_horiz_address_in_valid 	),
	.horiz_address_in       (weight_1_horiz_address_in_bits		),
	.horiz_data_in_ready    (weight_1_horiz_data_in_ready    	),
	.horiz_data_in_valid    (weight_1_horiz_data_in_valid    	),
	.horiz_data_in          (weight_1_horiz_data_in_bits		),
	.PE_address_out_valid   (weight_1_PE_address_out_valid   	),
	.PE_address_out         (weight_1_PE_address_out_bits		),
	.PE_data_out_valid      (weight_1_PE_data_out_valid      	),
	.PE_data_out            (weight_1_PE_data_out_bits			),
	.horiz_address_out_ready(weight_1_horiz_address_out_ready	),
	.horiz_address_out_valid(weight_1_horiz_address_out_valid	),
	.horiz_address_out      (weight_1_horiz_address_out_bits	),
	.horiz_data_out_ready   (weight_1_horiz_data_out_ready   	),
	.horiz_data_out_valid   (weight_1_horiz_data_out_valid   	),
	.horiz_data_out         (weight_1_horiz_data_out_bits		),
	.data_in_sel            (weight_1_data_in_sel            	),
	.data_out_sel           (weight_1_data_out_sel           	)
);

Weight_Router Weight_Router_2 ( 
	.GLB_address_in_ready	(weight_2_GLB_address_in_ready	 	),
	.GLB_address_in_valid   (weight_2_GLB_address_in_valid   	),
	.GLB_address_in         (weight_2_GLB_address_in_bits		),
	.GLB_data_in_ready      (weight_2_GLB_data_in_ready      	),
	.GLB_data_in_valid      (weight_2_GLB_data_in_valid      	),
	.GLB_data_in            (weight_2_GLB_data_in_bits			),
	.horiz_address_in_ready (weight_2_horiz_address_in_ready 	),
	.horiz_address_in_valid (weight_2_horiz_address_in_valid 	),
	.horiz_address_in       (weight_2_horiz_address_in_bits		),
	.horiz_data_in_ready    (weight_2_horiz_data_in_ready    	),
	.horiz_data_in_valid    (weight_2_horiz_data_in_valid    	),
	.horiz_data_in          (weight_2_horiz_data_in_bits		),
	.PE_address_out_valid   (weight_2_PE_address_out_valid   	),
	.PE_address_out         (weight_2_PE_address_out_bits		),
	.PE_data_out_valid      (weight_2_PE_data_out_valid      	),
	.PE_data_out            (weight_2_PE_data_out_bits			),
	.horiz_address_out_ready(weight_2_horiz_address_out_ready	),
	.horiz_address_out_valid(weight_2_horiz_address_out_valid	),
	.horiz_address_out      (weight_2_horiz_address_out_bits	),
	.horiz_data_out_ready   (weight_2_horiz_data_out_ready   	),
	.horiz_data_out_valid   (weight_2_horiz_data_out_valid   	),
	.horiz_data_out         (weight_2_horiz_data_out_bits		),
	.data_in_sel            (weight_2_data_in_sel            	),
	.data_out_sel           (weight_2_data_out_sel           	)
);

Psum_Router Psum_Router_0 ( 
	.PE_in_ready    (psum_0_PE_in_ready    	),
	.PE_in_valid    (psum_0_PE_in_valid    	),
	.PE_in          (psum_0_PE_in_bits		),
	.GLB_in_ready   (psum_0_GLB_in_ready   	),
	.GLB_in_valid   (psum_0_GLB_in_valid   	),
	.GLB_in         (psum_0_GLB_in_bits		),
	.north_in_ready (psum_0_north_in_ready 	),
	.north_in_valid (psum_0_north_in_valid 	),
	.north_in       (psum_0_north_in_bits	),
	.PE_out_ready   (psum_0_PE_out_ready   	),
	.PE_out_valid   (psum_0_PE_out_valid   	),
	.PE_out         (psum_0_PE_out_bits		),
	.GLB_out_ready  (psum_0_GLB_out_ready  	),
	.GLB_out_valid  (psum_0_GLB_out_valid  	),
	.GLB_out		(psum_0_GLB_out_bits	),
	.south_out_ready(psum_0_south_out_ready	),
	.south_out_valid(psum_0_south_out_valid	),	
	.south_out      (psum_0_south_out_bits	),
	.data_in_sel    (psum_0_data_in_sel    	),
	.data_out_sel   (psum_0_data_out_sel   	)
);

Psum_Router Psum_Router_1 ( 
	.PE_in_ready    (psum_1_PE_in_ready    	),
	.PE_in_valid    (psum_1_PE_in_valid    	),
	.PE_in          (psum_1_PE_in_bits		),
	.GLB_in_ready   (psum_1_GLB_in_ready   	),
	.GLB_in_valid   (psum_1_GLB_in_valid   	),
	.GLB_in         (psum_1_GLB_in_bits		),
	.north_in_ready (psum_1_north_in_ready 	),
	.north_in_valid (psum_1_north_in_valid 	),
	.north_in       (psum_1_north_in_bits	),
	.PE_out_ready   (psum_1_PE_out_ready   	),
	.PE_out_valid   (psum_1_PE_out_valid   	),
	.PE_out         (psum_1_PE_out_bits		),
	.GLB_out_ready  (psum_1_GLB_out_ready  	),
	.GLB_out_valid  (psum_1_GLB_out_valid  	),
	.GLB_out		(psum_1_GLB_out_bits	),
	.south_out_ready(psum_1_south_out_ready	),
	.south_out_valid(psum_1_south_out_valid	),	
	.south_out      (psum_1_south_out_bits	),
	.data_in_sel    (psum_1_data_in_sel    	),
	.data_out_sel   (psum_1_data_out_sel   	)
);

Psum_Router Psum_Router_2 ( 
	.PE_in_ready    (psum_2_PE_in_ready    	),
	.PE_in_valid    (psum_2_PE_in_valid    	),
	.PE_in          (psum_2_PE_in_bits		),
	.GLB_in_ready   (psum_2_GLB_in_ready   	),
	.GLB_in_valid   (psum_2_GLB_in_valid   	),
	.GLB_in         (psum_2_GLB_in_bits		),
	.north_in_ready (psum_2_north_in_ready 	),
	.north_in_valid (psum_2_north_in_valid 	),
	.north_in       (psum_2_north_in_bits	),
	.PE_out_ready   (psum_2_PE_out_ready   	),
	.PE_out_valid   (psum_2_PE_out_valid   	),
	.PE_out         (psum_2_PE_out_bits		),
	.GLB_out_ready  (psum_2_GLB_out_ready  	),
	.GLB_out_valid  (psum_2_GLB_out_valid  	),
	.GLB_out		(psum_2_GLB_out_bits	),
	.south_out_ready(psum_2_south_out_ready	),
	.south_out_valid(psum_2_south_out_valid	),	
	.south_out      (psum_2_south_out_bits	),
	.data_in_sel    (psum_2_data_in_sel    	),
	.data_out_sel   (psum_2_data_out_sel   	)
);


endmodule
